`timescale 1ms/1ms

module main_t();


main mainTest();


endmodule
