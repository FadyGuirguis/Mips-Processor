module increment4(out, in);

input [9:0] in;
output [9:0] out;

assign out = in + 4;

endmodule